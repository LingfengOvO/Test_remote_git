'timescale 1ns\1ps
/***********************************************
#
#      Filename: test.v
#
#        Author: Clough - clough@gmail.com
#   Description: ---
#        Create: 2022-07-21 15:36:44
# Last Modified: 2022-07-22 14:48:47
***********************************************/

begin
    if( stream_out = 1'b1 ) begin
        
    end
    else if() begin

    end
end

begin
    
end
always @ (*)
begin
    if()
end
xiugai2
 
